// Copyright lowRISC contributors (OpenTitan project).
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

// Macro bodies included by prim_assert.sv for tools that support full SystemVerilog and SVA syntax.
// See prim_assert.sv for documentation for each of the macros.







































// NOTE: Removed default args for Quartus compatibility














// NOTE: Removed default args for Quartus compatibility






// NOTE: Removed default args for Quartus compatibility






// NOTE: Removed default args for Quartus compatibility





// NOTE: Removed default args for Quartus compatibility



 // NOTE: Removed default args for Quartus compatibility











