// Register with asynchronous reset.









///////////////////////////
// Macro for Sparse FSMs //
///////////////////////////






























